** sch_path: /home/timothyjabez/Documents/Open_Source_Circuit_Design/ISSCC_2025_V1/xschem/Benchmark_Circuits/test_analog/test_analog.sch
**.subckt test_analog
V6 vin_p GND 0.9 dc 0.9 ac 1 pulse(0 1 100p 100p 100p 1u 2u)
V7 vin_n GND 0.9
V8 VDD GND 1.8
V9 VSS GND 0
I0 VSS i_bias 10u
x1 VDD vout vin_p vin_n VSS i_bias en OpAmp
V1 en GND 1.8
C1 vout GND 1p m=1
**** begin user architecture code
.lib /usr/local/share/pdk/sky130B/libs.tech/combined/sky130.lib.spice tt
**** end user architecture code
**.ends

* expanding   symbol:  Benchmark_Circuits/OpAmp_Defect/OpAmp.sym # of pins=7
** sym_path: /home/timothyjabez/Documents/Open_Source_Circuit_Design/ISSCC_2025_V1/xschem/Benchmark_Circuits/OpAmp_Defect/OpAmp.sym
** sch_path: /home/timothyjabez/Documents/Open_Source_Circuit_Design/ISSCC_2025_V1/xschem/Benchmark_Circuits/OpAmp_Defect/OpAmp.sch
.subckt OpAmp VDD vout vin_p vin_n VSS i_bias en
*.ipin vin_p
*.ipin vin_n
*.iopin VSS
*.iopin VDD
*.opin vout
*.ipin i_bias
*.ipin en
XM1 vout Active_load_g VDD VDD sky130_fd_pr__pfet_01v8 L=1 W=8 nf=2 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM2 Active_load_g Active_load_g VDD VDD sky130_fd_pr__pfet_01v8 L=1 W=8 nf=2 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM3 Active_load_g vin_p I_mirror_d VSS sky130_fd_pr__nfet_01v8 L=0.5 W=16 nf=4 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM4 vout vin_n I_mirror_d VSS sky130_fd_pr__nfet_01v8 L=0.5 W=16 nf=4 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM5 I_mirror_d I_mirror_g VSS VSS sky130_fd_pr__nfet_01v8 L=1 W=8 nf=2 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=2 m=2
XM6 i_bias I_mirror_g VSS VSS sky130_fd_pr__nfet_01v8 L=1 W=8 nf=2 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM9 en_n en VDD VDD sky130_fd_pr__pfet_01v8 L=0.15 W=2 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM10 en_n en VSS VSS sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM7 i_bias en I_mirror_g VSS sky130_fd_pr__nfet_01v8 L=0.35 W=4 nf=2 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM8 I_mirror_g en_n VSS VSS sky130_fd_pr__nfet_01v8 L=0.35 W=4 nf=2 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM11 Active_load_g en VDD VDD sky130_fd_pr__pfet_01v8 L=0.35 W=4 nf=2 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
R_open R_open_p R_open_n 1G m=1
.ends

.GLOBAL GND
**** begin user architecture code




* ngspice commands
.options savecurrents

.control
save all

op
remzerovec

tran 100n 10u
plot v(vout)

meas tran trise_pulse TRIG v(vout) VAL=0.1*1.8 RISE=1 TARG v(vout) VAL=0.9*1.8 RISE=1
let slew_rate = 0.8*1.8/trise_pulse
print slew_rate > opamp_specs.txt
let power_consumption = -@V8[i]*v(VDD)
meas tran power_average AVG power_consumption from=0u to=10u
print power_average >> opamp_specs.txt
write top_level.out

set appendwrite
set units=degrees
dc V6 0 1.8 0.01
remzerovec
write top_level.out

ac dec 10 1 1e12
let gain = v(vout)/(v(vin_p)-v(vin_n))

; Measurement of OpAmp performance parameters
meas ac AOL_DC_dB FIND vdb(gain) AT=10 >> opamp_specs.txt
let gain_3dB = AOL_DC_dB-3
print gain_3dB
meas ac BW3dB when vdb(gain) = gain_3dB >> opamp_specs.txt
meas ac UGBW when vdb(gain) = 1 >> opamp_specs.txt
meas ac Phase_Unity_Gain FIND vp(gain) AT=UGBW >> opamp_specs.txt
meas ac Zero_PM_Freq when vp(gain)=-175 >> opamp_specs.txt
meas ac GM FIND vdb(gain) at=Zero_PM_Freq >> opamp_specs.txt
let PM = 180+Phase_Unity_Gain
print PM >> opamp_specs.txt

settype decibel gain
plot vdb(gain) ylabel 'gain mag'
plot cph(gain) ylabel 'gain phase'
write top_level.out
.endc


**** end user architecture code
.end
